package alu_pkg;

`include "alu_transaction.sv"
`include "alu_generator.sv"
`include "alu_driver_new.sv"
`include "alu_monitor.sv"
`include "reference_model_version1.sv"
`include "alu_scoreboard.sv"
`include "alu_environment.sv"
`include "alu_test.sv"

endpackage
